module plugboardEncode(input [4:0] code, output [4:0] val);	
	assign val = code;
endmodule
